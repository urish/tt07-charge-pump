* Dickson Charge Pump Teshbench

.include "pdk_lib.spice"

* Power supply
V1 VGND 0 0
V2 VPWR VGND 1.8
* Clock
V3 clk VGND PULSE(0 1.8 0 30p 30p {{PLACEHOLDER_CLOCK}})

* Load the output
R1 "ua[0]" 0 7.8Meg

.include "tt_um_urish_charge_pump.spice"

x1 clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
+ tt_um_urish_charge_pump

.tran 0.5n 50u

.control
run
wrdata voltage.txt "ua[0]"
.endc
.end

.end
